library verilog;
use verilog.vl_types.all;
entity CT2_vlg_vec_tst is
end CT2_vlg_vec_tst;
