library verilog;
use verilog.vl_types.all;
entity TRG_vlg_vec_tst is
end TRG_vlg_vec_tst;
