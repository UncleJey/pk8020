library verilog;
use verilog.vl_types.all;
entity Scheme_vlg_check_tst is
    port(
        out1_25         : in     vl_logic;
        out2_5          : in     vl_logic;
        out5            : in     vl_logic;
        out10           : in     vl_logic;
        out20           : in     vl_logic;
        out_LA2         : in     vl_logic;
        outC0           : in     vl_logic;
        outC1           : in     vl_logic;
        outC2           : in     vl_logic;
        outC3           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Scheme_vlg_check_tst;
