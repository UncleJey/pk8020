library verilog;
use verilog.vl_types.all;
entity T_vlg_vec_tst is
end T_vlg_vec_tst;
