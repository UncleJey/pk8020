library verilog;
use verilog.vl_types.all;
entity Scheme_vlg_vec_tst is
end Scheme_vlg_vec_tst;
